
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use WORK.VM2413.ALL;

entity VoiceRom is 
  port (  
    clk    : in std_logic;
    addr : in VOICE_ID_TYPE;
    data  : out VOICE_TYPE
  );
end VoiceRom;

architecture RTL of VoiceRom is

  type VOICE_ARRAY_TYPE is array (0 to 37) of VOICE_VECTOR_TYPE;
  constant voices : VOICE_ARRAY_TYPE := (
-- APEK<ML>KL< TL >W<F><AR><DR><SL><RR>
  "000000000000000000000000000000000000", -- @0(M)
  "000000000000000000000000000000000000", -- @0(C)
-- APEK<ML>KL< TL >W<F><AR><DR><SL><RR>
  "000000110000010101101110100001000010", -- @1(M)
  "001000010000000000001000000100100111", -- @1(C)
-- APEK<ML>KL< TL >W<F><AR><DR><SL><RR>
  "000100110001010011011101100000100011", -- @2(M)
  "010000010000000000001111011000010010", -- @2(C)
-- APEK<ML>KL< TL >W<F><AR><DR><SL><RR>
  "000100010000100010001111101000100000", -- @3(M)
  "000100010000000000001011001000010010", -- @3(C)
-- APEK<ML>KL< TL >W<F><AR><DR><SL><RR>
  "001100010000110001111010100001100001", -- @4(M)
  "011000010000000000000110010000100111", -- @4(C)
-- APEK<ML>KL< TL >W<F><AR><DR><SL><RR>
  "001100100001111001101110000100000001", -- @5(M)
  "001000010000000000000111011000101000", -- @5(C)
-- APEK<ML>KL< TL >W<F><AR><DR><SL><RR>
  "000000100000011000001010001111110100", -- @6(M)
  "000000010000000000001110001011110100", -- @6(C)
-- APEK<ML>KL< TL >W<F><AR><DR><SL><RR>
  "001000010001110101111000001000010001", -- @7(M)
  "011000010000000000001000000100000111", -- @7(C)
-- APEK<ML>KL< TL >W<F><AR><DR><SL><RR>
  "001000110010001001111010001000000001", -- @8(M)
  "001000010000000010000111001000010111", -- @8(C)
-- APEK<ML>KL< TL >W<F><AR><DR><SL><RR>
  "001101010010010100000100000001110010", -- @9(M)
  "000100010000000000000111001100000001", -- @9(C)
-- APEK<ML>KL< TL >W<F><AR><DR><SL><RR>
  "101101010000111111111010100001010001", -- @10(M)
  "000000010000000000001010010100000010", -- @10(C)
-- APEK<ML>KL< TL >W<F><AR><DR><SL><RR>
  "000101110010010001111111100000100010", -- @11(M)
  "110000010000000000001111100000010010", -- @11(C)
-- APEK<ML>KL< TL >W<F><AR><DR><SL><RR>
  "011100010001000101100110010100011000", -- @12(M)
  "001000110000000000000111010000010110", -- @12(C)
-- APEK<ML>KL< TL >W<F><AR><DR><SL><RR>
  "000000011101001101011100100100000011", -- @13(M)
  "000000100000000000001001010100000010", -- @13(C)
-- APEK<ML>KL< TL >W<F><AR><DR><SL><RR>
  "011000010000110000001001010000110011", -- @14(M)
  "011000110000000000001100000011110110", -- @14(C)
-- APEK<ML>KL< TL >W<F><AR><DR><SL><RR>
  "001000010000110100001100000101010110", -- @15(M)
  "011100100000000000001101010100000110", -- @15(C)
-- APEK<ML>KL< TL >W<F><AR><DR><SL><RR>
  "000000010001100011111101111101101010", -- @16(M)
  "000000010000000000001111100001101101", -- @16(C)
-- APEK<ML>KL< TL >W<F><AR><DR><SL><RR>
  "000000010000000000001100100010100111", -- @17(M)
  "000000010000000000001101100001101000", -- @17(C)
-- APEK<ML>KL< TL >W<F><AR><DR><SL><RR>
  "000001010000000000001111100001011001", -- @18(M)
  "000000010000000000001010101001010101"  -- @18(C)
);

begin

  process (clk) 

  begin
  
    if clk'event and clk = '1' then
	  data <= CONV_VOICE(voices(addr));
    end if;
    
  end process;

end RTL;