
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use WORK.VM2413.ALL;

entity VoiceRom is 
  port (  
    clk    : in std_logic;
    addr : in VOICE_ID_TYPE;
    data  : out VOICE_TYPE
  );
end VoiceRom;

architecture RTL of VoiceRom is

  type VOICE_ARRAY_TYPE is array (0 to 37) of VOICE_VECTOR_TYPE;
  constant voices : VOICE_ARRAY_TYPE := (
-- APEK<ML>KL< TL >W<F><AR><DR><SL><RR>
  "000000000000000000000000000000000000", -- @0(M)
  "000000000000000000000000000000000000", -- @0(C)
-- APEK<ML>KL< TL >W<F><AR><DR><SL><RR>
  "001100110000100111101001010001000000", -- @1(M)
  "000000010000000000001001000000000001", -- @1(C)
-- APEK<ML>KL< TL >W<F><AR><DR><SL><RR>
  "000100110000111111011100111001000011", -- @2(M)
  "010000010000000000001101001100010011", -- @2(C)
-- APEK<ML>KL< TL >W<F><AR><DR><SL><RR>
  "000000010001101101101111111100000000", -- @3(M)
  "000100100000000000001101001000110010", -- @3(C)
-- APEK<ML>KL< TL >W<F><AR><DR><SL><RR>
  "011000010001101101111010111100100000", -- @4(M)
  "011000010000000000000110001100101000", -- @4(C)
-- APEK<ML>KL< TL >W<F><AR><DR><SL><RR>
  "001000100001111001101111000000001000", -- @5(M)
  "001000010000000000000111011000101000", -- @5(C)
-- APEK<ML>KL< TL >W<F><AR><DR><SL><RR>
  "011001100001010100001001001100100000", -- @6(M)
  "001000010000000000001001010011111000", -- @6(C)
-- APEK<ML>KL< TL >W<F><AR><DR><SL><RR>
  "001000010001110001111000001000010000", -- @7(M)
  "011000010000000000001000000100010111", -- @7(C)
-- APEK<ML>KL< TL >W<F><AR><DR><SL><RR>
  "001000110010000011111100000000000111", -- @8(M)
  "001000010000000010000111000101000111", -- @8(C)
-- APEK<ML>KL< TL >W<F><AR><DR><SL><RR>
  "001001010010011001010110010000011000", -- @9(M)
  "001100010000000000000100000111111000", -- @9(C)
-- APEK<ML>KL< TL >W<F><AR><DR><SL><RR>
  "000101110010100001111111111100000010", -- @10(M)
  "001000010000000000001000001111111000", -- @10(C)
-- APEK<ML>KL< TL >W<F><AR><DR><SL><RR>
  "100101110010010101111100111100000010", -- @11(M)
  "100000010000000000001100100000010100", -- @11(C)
-- APEK<ML>KL< TL >W<F><AR><DR><SL><RR>
  "001000010101010011111000000000000111", -- @12(M)
  "001000010000000000000111111100000111", -- @12(C)
-- APEK<ML>KL< TL >W<F><AR><DR><SL><RR>
  "000000010101011000111101001101000011", -- @13(M)
  "000000010000000000001011001001011000", -- @13(C)
-- APEK<ML>KL< TL >W<F><AR><DR><SL><RR>
  "001100010000110000111000001001000000", -- @14(M)
  "001000010000000000001100000000000111", -- @14(C)
-- APEK<ML>KL< TL >W<F><AR><DR><SL><RR>
  "001000010000110000111101010001000000", -- @15(M)
  "000000010000000000001101001110000100", -- @15(C)
-- APEK<ML>KL< TL >W<F><AR><DR><SL><RR>
  "000001000010100000001101111111111111", -- @16(M)
  "001000010000000000001111100011111000", -- @16(C)
-- APEK<ML>KL< TL >W<F><AR><DR><SL><RR>
  "001000110000000000001010100011111000", -- @17(M)
  "001000100000000000001111100011111000", -- @17(C)
-- APEK<ML>KL< TL >W<F><AR><DR><SL><RR>
  "001001010000000000001111100011111000", -- @18(M)
  "000110000000000000001010100101010101" -- @18(C)
);

begin

  process (clk) 

  begin
  
    if clk'event and clk = '1' then
	  data <= CONV_VOICE(voices(addr));
    end if;
    
  end process;

end RTL;